*******************************************************************************
* CDL netlist
*
* Library : LibreriaBruschi
* Top Cell Name: OTAPMOS
* View Name: extracted
* Netlist created: 23.lug.2019 18:29:34
*******************************************************************************

*.SCALE METER
*.GLOBAL 

*******************************************************************************
* Library Name: LibreriaBruschi
* Cell Name:    OTAPMOS
* View Name:    extracted
*******************************************************************************

.SUBCKT OTAPMOS

MM39 n1 n8 n0 n0 N_PSM025 w=6e-06 l=1e-06 as=7.5e-12 ps=1.45e-05 ad=7.5e-12 pd=1.45e-05 $X=59.6 $Y=4.1
MM43 n7 n8 n0 n0 N_PSM025 w=6e-06 l=1e-06 as=7.5e-12 ps=1.45e-05 ad=7.5e-12 pd=1.45e-05 $X=128.65 $Y=4.1
MM50 n2 n1 n1 n2 P_PSM025 w=2.6e-05 l=1e-06 as=3.12e-11 ps=5.44e-05 ad=2.86e-11 pd=5.42e-05 $X=103.8 $Y=24.5
MM41 n3 n3 n0 n0 N_PSM025 w=6e-06 l=1e-06 as=7.5e-12 ps=1.45e-05 ad=7.5e-12 pd=1.45e-05 $X=87.15 $Y=4.1
MM47 n6 n9 n8 n2 P_PSM025 w=1.3e-05 l=1e-06 as=1.3e-11 ps=2.8e-05 ad=1.3e-11 pd=2.8e-05 $X=64.05 $Y=14.75
MM51 n2 n1 n4 n2 P_PSM025 w=2.6e-05 l=1e-06 as=3.12e-11 ps=5.44e-05 ad=2.86e-11 pd=5.42e-05 $X=134.55 $Y=24.5
MM42 n4 n3 n0 n0 N_PSM025 w=6e-06 l=1e-06 as=7.5e-12 ps=1.45e-05 ad=7.5e-12 pd=1.45e-05 $X=96 $Y=4.1
MM44 n7 n3 n0 n0 N_PSM025 w=6e-06 l=1e-06 as=7.5e-12 ps=1.45e-05 ad=7.5e-12 pd=1.45e-05 $X=139 $Y=4.1
MM45 n2 n4 n7 n0 N_PSM025 w=1.2e-05 l=1e-06 as=1.86e-11 ps=2.71e-05 ad=1.74e-11 pd=2.69e-05 $X=150.6 $Y=4
MM48 n2 n5 n6 n2 P_PSM025 w=2.6e-05 l=1e-06 as=3.12e-11 ps=5.44e-05 ad=2.86e-11 pd=5.42e-05 $X=73.3 $Y=24.5
MM40 n8 n8 n0 n0 N_PSM025 w=6e-06 l=1e-06 as=7.5e-12 ps=1.45e-05 ad=7.5e-12 pd=1.45e-05 $X=67.75 $Y=4.1
MM49 n6 n10 n3 n2 P_PSM025 w=1.3e-05 l=1e-06 as=1.3e-11 ps=2.8e-05 ad=1.3e-11 pd=2.8e-05 $X=83.1 $Y=14.75
MM46 n2 n5 n5 n2 P_PSM025 w=2.6e-05 l=1e-06 as=3.12e-11 ps=5.44e-05 ad=2.86e-11 pd=5.42e-05 $X=44.15 $Y=24.5
.ENDS
